module terminal_top(
  input clk,
  input resetn,

  output       tmds_clk_n,
  output       tmds_clk_p,
  output [2:0] tmds_d_n,
  output [2:0] tmds_d_p
);

  clock_generator clk_gen (
    .clkout(clk_p5), //output clkout
    .lock(pll_lock), //output lock
    .clkin(clk) //input clkin
  );

  clock_div5 clk_div (
    .clkout(clk_p), //output clkout
    .hclkin(clk_p5), //input hclkin
    .resetn(pll_lock) //input resetn
  );

  hdmi_term terminal (
    .clk(clk_p),
    .resetn(sys_resetn),

    // video clocks
    .clk_pixel(clk_p),
    .clk_5x_pixel(clk_p5),
    .locked(pll_lock),

    // output signals
    .tmds_clk_n(tmds_clk_n),
    .tmds_clk_p(tmds_clk_p),
    .tmds_d_n(tmds_d_n),
    .tmds_d_p(tmds_d_p)
  );

  Reset_Sync u_Reset_Sync (
    .resetn(sys_resetn),
    .ext_reset(resetn & pll_lock),
    .clk(clk_p)
  );

endmodule

module Reset_Sync (
 input clk,
 input ext_reset,
 output resetn
);

 reg [3:0] reset_cnt = 0;
 
 always @(posedge clk or negedge ext_reset) begin
     if (~ext_reset)
         reset_cnt <= 4'b0;
     else
         reset_cnt <= reset_cnt + !resetn;
 end
 
 assign resetn = &reset_cnt;

endmodule